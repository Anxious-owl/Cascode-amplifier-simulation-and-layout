magic
tech scmos
timestamp 1731230711
<< nwell >>
rect -34 0 120 66
<< ntransistor >>
rect -16 -22 -14 -17
rect 22 -27 24 -17
rect 60 -27 62 -17
rect 98 -27 100 -17
rect 6 -57 8 -47
rect 42 -57 44 -47
rect 78 -57 80 -47
<< ptransistor >>
rect -20 15 -18 39
rect 10 15 12 39
rect 41 31 43 39
rect 73 15 75 39
rect 104 15 106 39
<< ndiffusion >>
rect -20 -22 -16 -17
rect -14 -22 -10 -17
rect 18 -27 22 -17
rect 24 -27 28 -17
rect 56 -27 60 -17
rect 62 -27 66 -17
rect 94 -27 98 -17
rect 100 -27 104 -17
rect 2 -57 6 -47
rect 8 -57 12 -47
rect 38 -57 42 -47
rect 44 -57 48 -47
rect 74 -57 78 -47
rect 80 -57 84 -47
<< pdiffusion >>
rect -24 34 -20 39
rect -28 29 -20 34
rect -24 24 -20 29
rect -28 20 -20 24
rect -24 15 -20 20
rect -18 15 -14 39
rect 6 34 10 39
rect 2 29 10 34
rect 6 24 10 29
rect 2 20 10 24
rect 6 15 10 20
rect 12 34 16 39
rect 12 29 20 34
rect 36 31 41 39
rect 43 31 48 39
rect 68 34 73 39
rect 12 24 16 29
rect 64 29 73 34
rect 12 20 20 24
rect 12 15 16 20
rect 68 24 73 29
rect 64 20 73 24
rect 68 15 73 20
rect 75 34 80 39
rect 75 29 84 34
rect 75 24 80 29
rect 75 20 84 24
rect 75 15 80 20
rect 100 34 104 39
rect 96 29 104 34
rect 100 24 104 29
rect 96 20 104 24
rect 100 15 104 20
rect 106 34 110 39
rect 106 29 114 34
rect 106 24 110 29
rect 106 20 114 24
rect 106 15 110 20
<< ndcontact >>
rect -24 -22 -20 -17
rect -10 -22 -6 -17
rect 14 -27 18 -17
rect 28 -27 32 -17
rect 52 -27 56 -17
rect 66 -27 70 -17
rect 90 -27 94 -17
rect 104 -27 108 -17
rect -2 -57 2 -47
rect 12 -57 16 -47
rect 34 -57 38 -47
rect 48 -57 52 -47
rect 70 -57 74 -47
rect 84 -57 88 -47
<< pdcontact >>
rect -28 34 -24 39
rect -28 24 -24 29
rect -28 15 -24 20
rect -14 15 -10 39
rect 2 34 6 39
rect 2 24 6 29
rect 2 15 6 20
rect 16 34 20 39
rect 32 31 36 39
rect 48 31 52 39
rect 64 34 68 39
rect 16 24 20 29
rect 16 15 20 20
rect 64 24 68 29
rect 64 15 68 20
rect 80 34 84 39
rect 80 24 84 29
rect 80 15 84 20
rect 96 34 100 39
rect 96 24 100 29
rect 96 15 100 20
rect 110 34 114 39
rect 110 24 114 29
rect 110 15 114 20
<< psubstratepcontact >>
rect -20 -73 -15 -67
rect 9 -73 14 -67
rect 45 -73 50 -67
rect 75 -73 80 -67
rect 102 -73 107 -67
<< nsubstratencontact >>
rect -24 56 -19 62
rect 6 56 11 62
rect 36 56 41 62
rect 68 56 73 62
rect 100 56 105 62
<< polysilicon >>
rect -20 39 -18 43
rect 10 39 12 43
rect 41 39 43 43
rect 73 39 75 43
rect 104 39 106 43
rect 41 30 43 31
rect -20 13 -18 15
rect 10 13 12 15
rect 73 13 75 15
rect 104 14 106 15
rect -16 -17 -14 -14
rect 22 -17 24 -14
rect 60 -17 62 -14
rect 98 -17 100 -13
rect -16 -27 -14 -22
rect 22 -33 24 -27
rect 60 -30 62 -27
rect 98 -33 100 -27
rect 6 -47 8 -44
rect 42 -47 44 -44
rect 78 -47 80 -44
rect 6 -59 8 -57
rect 42 -59 44 -57
rect 78 -59 80 -57
<< polycontact >>
rect 40 26 44 30
rect -21 8 -17 13
rect 9 8 13 13
rect 72 9 76 13
rect 103 10 107 14
rect -17 -14 -13 -10
rect 21 -14 25 -10
rect 59 -14 63 -10
rect 97 -13 101 -9
rect -17 -31 -13 -27
rect 59 -34 63 -30
rect 5 -63 9 -59
rect 41 -63 45 -59
rect 77 -63 81 -59
<< metal1 >>
rect -30 56 -24 62
rect -19 56 6 62
rect 11 56 36 62
rect 41 56 68 62
rect 73 56 100 62
rect 105 56 117 62
rect -28 39 -24 56
rect 2 39 6 56
rect 32 39 36 56
rect 64 48 91 52
rect 64 39 68 48
rect -28 29 -24 34
rect -28 20 -24 24
rect 2 29 6 34
rect 64 29 68 34
rect 2 20 6 24
rect 64 20 68 24
rect -26 9 -21 12
rect -17 9 9 12
rect 88 6 91 48
rect 96 39 100 56
rect 96 29 100 34
rect 96 20 100 24
rect 110 29 114 34
rect 110 20 114 24
rect 110 6 114 15
rect 88 3 114 6
rect -13 -13 21 -10
rect -10 -17 -6 -13
rect 25 -13 59 -10
rect 63 -13 97 -10
rect -24 -73 -20 -22
rect 14 -33 18 -27
rect 52 -33 56 -27
rect 12 -37 18 -33
rect 48 -37 56 -33
rect 90 -33 94 -27
rect 84 -37 94 -33
rect 12 -47 16 -37
rect 48 -47 52 -37
rect 84 -47 88 -37
rect -2 -67 2 -57
rect 34 -67 38 -57
rect 70 -67 74 -57
rect -15 -73 9 -67
rect 14 -73 45 -67
rect 50 -73 75 -67
rect 80 -73 102 -67
rect 107 -73 111 -67
<< metal2 >>
rect -14 -1 -10 39
rect 16 -1 20 39
rect 40 23 44 30
rect 48 23 52 39
rect 40 20 52 23
rect 40 13 44 20
rect 80 14 84 39
rect 40 9 76 13
rect 40 -1 44 9
rect 72 6 76 9
rect 80 11 121 14
rect 80 -1 84 11
rect -14 -5 5 -1
rect 16 -5 32 -1
rect 40 -5 70 -1
rect 1 -27 5 -5
rect -17 -31 5 -27
rect 28 -59 32 -5
rect 66 -27 70 -5
rect 80 -6 108 -1
rect 104 -27 108 -6
rect 59 -37 63 -33
rect 5 -62 84 -59
<< labels >>
rlabel metal1 42 59 42 59 1 vdd!
rlabel metal1 43 -70 43 -70 1 gnd!
rlabel metal1 -24 10 -24 10 1 vbiasp
rlabel metal1 44 -11 44 -11 1 vbias3
rlabel metal2 106 -4 106 -4 1 vbias1
rlabel metal2 68 -4 68 -4 1 vbias2
rlabel metal2 30 -35 30 -35 1 vbias4
rlabel metal2 -12 -2 -12 -2 1 test1
<< end >>
